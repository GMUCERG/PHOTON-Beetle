
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;


entity mcs_rom is
	generic(sel : integer := 0);
	port(ADDR : in  STD_LOGIC_VECTOR(4 downto 0);
	     Dout : out STD_LOGIC_VECTOR(3 downto 0));
end mcs_rom;

architecture mr0 of mcs_rom is

	signal input1 : integer range 0 to 31;
	type v_arr is array (0 to 31) of STD_LOGIC_VECTOR(3 downto 0);

begin

	gen_mcs_rom : -- Cell 0 :: 2 | 2 --
	if sel = 0 generate
		constant MEMORY : v_arr := ("0000",
		                            "0010",
		                            "0100",
		                            "0110",
		                            "1000",
		                            "1010",
		                            "1100",
		                            "1110",
		                            "0011",
		                            "0001",
		                            "0111",
		                            "0101",
		                            "1011",
		                            "1001",
		                            "1111",
		                            "1101",
		                            "0000",
		                            "0010",
		                            "0100",
		                            "0110",
		                            "1000",
		                            "1010",
		                            "1100",
		                            "1110",
		                            "0011",
		                            "0001",
		                            "0111",
		                            "0101",
		                            "1011",
		                            "1001",
		                            "1111",
		                            "1101");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 1 :: 4 | 8 --
	end generate;
    gen_mcs_rom_1: if sel = 1 generate

		constant MEMORY : v_arr := ("0000",
		                            "0100",
		                            "1000",
		                            "1100",
		                            "0011",
		                            "0111",
		                            "1011",
		                            "1111",
		                            "0110",
		                            "0010",
		                            "1110",
		                            "1010",
		                            "0101",
		                            "0001",
		                            "1101",
		                            "1001",
		                            "0000",
		                            "1000",
		                            "0011",
		                            "1011",
		                            "0110",
		                            "1110",
		                            "0101",
		                            "1101",
		                            "1100",
		                            "0100",
		                            "1111",
		                            "0111",
		                            "1010",
		                            "0010",
		                            "1001",
		                            "0001");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 2 :: 2 | 5 --
	end generate;
    gen_mcs_rom_2: if sel = 2 generate

		constant MEMORY : v_arr := ("0000",
		                            "0010",
		                            "0100",
		                            "0110",
		                            "1000",
		                            "1010",
		                            "1100",
		                            "1110",
		                            "0011",
		                            "0001",
		                            "0111",
		                            "0101",
		                            "1011",
		                            "1001",
		                            "1111",
		                            "1101",
		                            "0000",
		                            "0101",
		                            "1010",
		                            "1111",
		                            "0111",
		                            "0010",
		                            "1101",
		                            "1000",
		                            "1110",
		                            "1011",
		                            "0100",
		                            "0001",
		                            "1001",
		                            "1100",
		                            "0011",
		                            "0110");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 3 :: 11 | 6 --
	end generate;
    gen_mcs_rom_3: if sel = 3 generate

		constant MEMORY : v_arr := ("0000",
		                            "1011",
		                            "0101",
		                            "1110",
		                            "1010",
		                            "0001",
		                            "1111",
		                            "0100",
		                            "0111",
		                            "1100",
		                            "0010",
		                            "1001",
		                            "1101",
		                            "0110",
		                            "1000",
		                            "0011",
		                            "0000",
		                            "0110",
		                            "1100",
		                            "1010",
		                            "1011",
		                            "1101",
		                            "0111",
		                            "0001",
		                            "0101",
		                            "0011",
		                            "1001",
		                            "1111",
		                            "1110",
		                            "1000",
		                            "0010",
		                            "0100");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 4 :: 12 | 7 --
	end generate;
    gen_mcs_rom_4: if sel = 4 generate

		constant MEMORY : v_arr := ("0000",
		                            "1100",
		                            "1011",
		                            "0111",
		                            "0101",
		                            "1001",
		                            "1110",
		                            "0010",
		                            "1010",
		                            "0110",
		                            "0001",
		                            "1101",
		                            "1111",
		                            "0011",
		                            "0100",
		                            "1000",
		                            "0000",
		                            "0111",
		                            "1110",
		                            "1001",
		                            "1111",
		                            "1000",
		                            "0001",
		                            "0110",
		                            "1101",
		                            "1010",
		                            "0011",
		                            "0100",
		                            "0010",
		                            "0101",
		                            "1100",
		                            "1011");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 5 :: 9 | 7 --
	end generate;
    gen_mcs_rom_5: if sel = 5 generate

		constant MEMORY : v_arr := ("0000",
		                            "1001",
		                            "0001",
		                            "1000",
		                            "0010",
		                            "1011",
		                            "0011",
		                            "1010",
		                            "0100",
		                            "1101",
		                            "0101",
		                            "1100",
		                            "0110",
		                            "1111",
		                            "0111",
		                            "1110",
		                            "0000",
		                            "0111",
		                            "1110",
		                            "1001",
		                            "1111",
		                            "1000",
		                            "0001",
		                            "0110",
		                            "1101",
		                            "1010",
		                            "0011",
		                            "0100",
		                            "0010",
		                            "0101",
		                            "1100",
		                            "1011");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 6 :: 8 | 5 --
	end generate;
    gen_mcs_rom_6: if sel = 6 generate

		constant MEMORY : v_arr := ("0000",
		                            "1000",
		                            "0011",
		                            "1011",
		                            "0110",
		                            "1110",
		                            "0101",
		                            "1101",
		                            "1100",
		                            "0100",
		                            "1111",
		                            "0111",
		                            "1010",
		                            "0010",
		                            "1001",
		                            "0001",
		                            "0000",
		                            "0101",
		                            "1010",
		                            "1111",
		                            "0111",
		                            "0010",
		                            "1101",
		                            "1000",
		                            "1110",
		                            "1011",
		                            "0100",
		                            "0001",
		                            "1001",
		                            "1100",
		                            "0011",
		                            "0110");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 7 :: 13 | 2 --
	end generate;
    gen_mcs_rom_7: if sel = 7 generate

		constant MEMORY : v_arr := ("0000",
		                            "1101",
		                            "1001",
		                            "0100",
		                            "0001",
		                            "1100",
		                            "1000",
		                            "0101",
		                            "0010",
		                            "1111",
		                            "1011",
		                            "0110",
		                            "0011",
		                            "1110",
		                            "1010",
		                            "0111",
		                            "0000",
		                            "0010",
		                            "0100",
		                            "0110",
		                            "1000",
		                            "1010",
		                            "1100",
		                            "1110",
		                            "0011",
		                            "0001",
		                            "0111",
		                            "0101",
		                            "1011",
		                            "1001",
		                            "1111",
		                            "1101");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 8 :: 4 | 9 --
	end generate;
    gen_mcs_rom_8: if sel = 8 generate

		constant MEMORY : v_arr := ("0000",
		                            "0100",
		                            "1000",
		                            "1100",
		                            "0011",
		                            "0111",
		                            "1011",
		                            "1111",
		                            "0110",
		                            "0010",
		                            "1110",
		                            "1010",
		                            "0101",
		                            "0001",
		                            "1101",
		                            "1001",
		                            "0000",
		                            "1001",
		                            "0001",
		                            "1000",
		                            "0010",
		                            "1011",
		                            "0011",
		                            "1010",
		                            "0100",
		                            "1101",
		                            "0101",
		                            "1100",
		                            "0110",
		                            "1111",
		                            "0111",
		                            "1110");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 9 :: 4 | 4 --
	end generate;
    gen_mcs_rom_9: if sel = 9 generate

		constant MEMORY : v_arr := ("0000",
		                            "0100",
		                            "1000",
		                            "1100",
		                            "0011",
		                            "0111",
		                            "1011",
		                            "1111",
		                            "0110",
		                            "0010",
		                            "1110",
		                            "1010",
		                            "0101",
		                            "0001",
		                            "1101",
		                            "1001",
		                            "0000",
		                            "0100",
		                            "1000",
		                            "1100",
		                            "0011",
		                            "0111",
		                            "1011",
		                            "1111",
		                            "0110",
		                            "0010",
		                            "1110",
		                            "1010",
		                            "0101",
		                            "0001",
		                            "1101",
		                            "1001");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 10 :: 13 | 13 --
	end generate;
    gen_mcs_rom_10: if sel = 10 generate

		constant MEMORY : v_arr := ("0000",
		                            "1101",
		                            "1001",
		                            "0100",
		                            "0001",
		                            "1100",
		                            "1000",
		                            "0101",
		                            "0010",
		                            "1111",
		                            "1011",
		                            "0110",
		                            "0011",
		                            "1110",
		                            "1010",
		                            "0111",
		                            "0000",
		                            "1101",
		                            "1001",
		                            "0100",
		                            "0001",
		                            "1100",
		                            "1000",
		                            "0101",
		                            "0010",
		                            "1111",
		                            "1011",
		                            "0110",
		                            "0011",
		                            "1110",
		                            "1010",
		                            "0111");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 11 :: 13 | 9 --
	end generate;
    gen_mcs_rom_11: if sel = 11 generate

		constant MEMORY : v_arr := ("0000",
		                            "1101",
		                            "1001",
		                            "0100",
		                            "0001",
		                            "1100",
		                            "1000",
		                            "0101",
		                            "0010",
		                            "1111",
		                            "1011",
		                            "0110",
		                            "0011",
		                            "1110",
		                            "1010",
		                            "0111",
		                            "0000",
		                            "1001",
		                            "0001",
		                            "1000",
		                            "0010",
		                            "1011",
		                            "0011",
		                            "1010",
		                            "0100",
		                            "1101",
		                            "0101",
		                            "1100",
		                            "0110",
		                            "1111",
		                            "0111",
		                            "1110");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 12 :: 1 | 12 --
	end generate;
    gen_mcs_rom_12: if sel = 12 generate

		constant MEMORY : v_arr := ("0000",
		                            "0001",
		                            "0010",
		                            "0011",
		                            "0100",
		                            "0101",
		                            "0110",
		                            "0111",
		                            "1000",
		                            "1001",
		                            "1010",
		                            "1011",
		                            "1100",
		                            "1101",
		                            "1110",
		                            "1111",
		                            "0000",
		                            "1100",
		                            "1011",
		                            "0111",
		                            "0101",
		                            "1001",
		                            "1110",
		                            "0010",
		                            "1010",
		                            "0110",
		                            "0001",
		                            "1101",
		                            "1111",
		                            "0011",
		                            "0100",
		                            "1000");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 13 :: 6 | 13 --
	end generate;
    gen_mcs_rom_13: if sel = 13 generate

		constant MEMORY : v_arr := ("0000",
		                            "0110",
		                            "1100",
		                            "1010",
		                            "1011",
		                            "1101",
		                            "0111",
		                            "0001",
		                            "0101",
		                            "0011",
		                            "1001",
		                            "1111",
		                            "1110",
		                            "1000",
		                            "0010",
		                            "0100",
		                            "0000",
		                            "1101",
		                            "1001",
		                            "0100",
		                            "0001",
		                            "1100",
		                            "1000",
		                            "0101",
		                            "0010",
		                            "1111",
		                            "1011",
		                            "0110",
		                            "0011",
		                            "1110",
		                            "1010",
		                            "0111");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 14 :: 5 | 15 --
	end generate;
    gen_mcs_rom_14: if sel = 14 generate

		constant MEMORY : v_arr := ("0000",
		                            "0101",
		                            "1010",
		                            "1111",
		                            "0111",
		                            "0010",
		                            "1101",
		                            "1000",
		                            "1110",
		                            "1011",
		                            "0100",
		                            "0001",
		                            "1001",
		                            "1100",
		                            "0011",
		                            "0110",
		                            "0000",
		                            "1111",
		                            "1101",
		                            "0010",
		                            "1001",
		                            "0110",
		                            "0100",
		                            "1011",
		                            "0001",
		                            "1110",
		                            "1100",
		                            "0011",
		                            "1000",
		                            "0111",
		                            "0101",
		                            "1010");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 15 :: 1 | 14 --
	end generate;
    gen_mcs_rom_15: if sel = 15 generate

		constant MEMORY : v_arr := ("0000",
		                            "0001",
		                            "0010",
		                            "0011",
		                            "0100",
		                            "0101",
		                            "0110",
		                            "0111",
		                            "1000",
		                            "1001",
		                            "1010",
		                            "1011",
		                            "1100",
		                            "1101",
		                            "1110",
		                            "1111",
		                            "0000",
		                            "1110",
		                            "1111",
		                            "0001",
		                            "1101",
		                            "0011",
		                            "0010",
		                            "1100",
		                            "1001",
		                            "0111",
		                            "0110",
		                            "1000",
		                            "0100",
		                            "1010",
		                            "1011",
		                            "0101");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 16 :: 15 | 14 --
	end generate;
    gen_mcs_rom_16: if sel = 16 generate

		constant MEMORY : v_arr := ("0000",
		                            "1111",
		                            "1101",
		                            "0010",
		                            "1001",
		                            "0110",
		                            "0100",
		                            "1011",
		                            "0001",
		                            "1110",
		                            "1100",
		                            "0011",
		                            "1000",
		                            "0111",
		                            "0101",
		                            "1010",
		                            "0000",
		                            "1110",
		                            "1111",
		                            "0001",
		                            "1101",
		                            "0011",
		                            "0010",
		                            "1100",
		                            "1001",
		                            "0111",
		                            "0110",
		                            "1000",
		                            "0100",
		                            "1010",
		                            "1011",
		                            "0101");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 17 :: 12 | 5 --
	end generate;
    gen_mcs_rom_17: if sel = 17 generate

		constant MEMORY : v_arr := ("0000",
		                            "1100",
		                            "1011",
		                            "0111",
		                            "0101",
		                            "1001",
		                            "1110",
		                            "0010",
		                            "1010",
		                            "0110",
		                            "0001",
		                            "1101",
		                            "1111",
		                            "0011",
		                            "0100",
		                            "1000",
		                            "0000",
		                            "0101",
		                            "1010",
		                            "1111",
		                            "0111",
		                            "0010",
		                            "1101",
		                            "1000",
		                            "1110",
		                            "1011",
		                            "0100",
		                            "0001",
		                            "1001",
		                            "1100",
		                            "0011",
		                            "0110");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 18 :: 9 | 14 --
	end generate;
    gen_mcs_rom_18: if sel = 18 generate

		constant MEMORY : v_arr := ("0000",
		                            "1001",
		                            "0001",
		                            "1000",
		                            "0010",
		                            "1011",
		                            "0011",
		                            "1010",
		                            "0100",
		                            "1101",
		                            "0101",
		                            "1100",
		                            "0110",
		                            "1111",
		                            "0111",
		                            "1110",
		                            "0000",
		                            "1110",
		                            "1111",
		                            "0001",
		                            "1101",
		                            "0011",
		                            "0010",
		                            "1100",
		                            "1001",
		                            "0111",
		                            "0110",
		                            "1000",
		                            "0100",
		                            "1010",
		                            "1011",
		                            "0101");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 19 :: 13 | 13 --
	end generate;
    gen_mcs_rom_19: if sel = 19 generate

		constant MEMORY : v_arr := ("0000",
		                            "1101",
		                            "1001",
		                            "0100",
		                            "0001",
		                            "1100",
		                            "1000",
		                            "0101",
		                            "0010",
		                            "1111",
		                            "1011",
		                            "0110",
		                            "0011",
		                            "1110",
		                            "1010",
		                            "0111",
		                            "0000",
		                            "1101",
		                            "1001",
		                            "0100",
		                            "0001",
		                            "1100",
		                            "1000",
		                            "0101",
		                            "0010",
		                            "1111",
		                            "1011",
		                            "0110",
		                            "0011",
		                            "1110",
		                            "1010",
		                            "0111");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 20 :: 9 | 4 --
	end generate;
    gen_mcs_rom_20: if sel = 20 generate

		constant MEMORY : v_arr := ("0000",
		                            "1001",
		                            "0001",
		                            "1000",
		                            "0010",
		                            "1011",
		                            "0011",
		                            "1010",
		                            "0100",
		                            "1101",
		                            "0101",
		                            "1100",
		                            "0110",
		                            "1111",
		                            "0111",
		                            "1110",
		                            "0000",
		                            "0100",
		                            "1000",
		                            "1100",
		                            "0011",
		                            "0111",
		                            "1011",
		                            "1111",
		                            "0110",
		                            "0010",
		                            "1110",
		                            "1010",
		                            "0101",
		                            "0001",
		                            "1101",
		                            "1001");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 21 :: 14 | 12 --
	end generate;
    gen_mcs_rom_21: if sel = 21 generate

		constant MEMORY : v_arr := ("0000",
		                            "1110",
		                            "1111",
		                            "0001",
		                            "1101",
		                            "0011",
		                            "0010",
		                            "1100",
		                            "1001",
		                            "0111",
		                            "0110",
		                            "1000",
		                            "0100",
		                            "1010",
		                            "1011",
		                            "0101",
		                            "0000",
		                            "1100",
		                            "1011",
		                            "0111",
		                            "0101",
		                            "1001",
		                            "1110",
		                            "0010",
		                            "1010",
		                            "0110",
		                            "0001",
		                            "1101",
		                            "1111",
		                            "0011",
		                            "0100",
		                            "1000");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 22 :: 5 | 9 --
	end generate;
    gen_mcs_rom_22: if sel = 22 generate

		constant MEMORY : v_arr := ("0000",
		                            "0101",
		                            "1010",
		                            "1111",
		                            "0111",
		                            "0010",
		                            "1101",
		                            "1000",
		                            "1110",
		                            "1011",
		                            "0100",
		                            "0001",
		                            "1001",
		                            "1100",
		                            "0011",
		                            "0110",
		                            "0000",
		                            "1001",
		                            "0001",
		                            "1000",
		                            "0010",
		                            "1011",
		                            "0011",
		                            "1010",
		                            "0100",
		                            "1101",
		                            "0101",
		                            "1100",
		                            "0110",
		                            "1111",
		                            "0111",
		                            "1110");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 23 :: 15 | 6 --
	end generate;
    gen_mcs_rom_23: if sel = 23 generate

		constant MEMORY : v_arr := ("0000",
		                            "1111",
		                            "1101",
		                            "0010",
		                            "1001",
		                            "0110",
		                            "0100",
		                            "1011",
		                            "0001",
		                            "1110",
		                            "1100",
		                            "0011",
		                            "1000",
		                            "0111",
		                            "0101",
		                            "1010",
		                            "0000",
		                            "0110",
		                            "1100",
		                            "1010",
		                            "1011",
		                            "1101",
		                            "0111",
		                            "0001",
		                            "0101",
		                            "0011",
		                            "1001",
		                            "1111",
		                            "1110",
		                            "1000",
		                            "0010",
		                            "0100");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 24 :: 12 | 3 --
	end generate;
    gen_mcs_rom_24: if sel = 24 generate

		constant MEMORY : v_arr := ("0000",
		                            "1100",
		                            "1011",
		                            "0111",
		                            "0101",
		                            "1001",
		                            "1110",
		                            "0010",
		                            "1010",
		                            "0110",
		                            "0001",
		                            "1101",
		                            "1111",
		                            "0011",
		                            "0100",
		                            "1000",
		                            "0000",
		                            "0011",
		                            "0110",
		                            "0101",
		                            "1100",
		                            "1111",
		                            "1010",
		                            "1001",
		                            "1011",
		                            "1000",
		                            "1101",
		                            "1110",
		                            "0111",
		                            "0100",
		                            "0001",
		                            "0010");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 25 :: 2 | 1 --
	end generate;
    gen_mcs_rom_25: if sel = 25 generate

		constant MEMORY : v_arr := ("0000",
		                            "0010",
		                            "0100",
		                            "0110",
		                            "1000",
		                            "1010",
		                            "1100",
		                            "1110",
		                            "0011",
		                            "0001",
		                            "0111",
		                            "0101",
		                            "1011",
		                            "1001",
		                            "1111",
		                            "1101",
		                            "0000",
		                            "0001",
		                            "0010",
		                            "0011",
		                            "0100",
		                            "0101",
		                            "0110",
		                            "0111",
		                            "1000",
		                            "1001",
		                            "1010",
		                            "1011",
		                            "1100",
		                            "1101",
		                            "1110",
		                            "1111");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 26 :: 2 | 1 --
	end generate;
    gen_mcs_rom_26: if sel = 26 generate

		constant MEMORY : v_arr := ("0000",
		                            "0010",
		                            "0100",
		                            "0110",
		                            "1000",
		                            "1010",
		                            "1100",
		                            "1110",
		                            "0011",
		                            "0001",
		                            "0111",
		                            "0101",
		                            "1011",
		                            "1001",
		                            "1111",
		                            "1101",
		                            "0000",
		                            "0001",
		                            "0010",
		                            "0011",
		                            "0100",
		                            "0101",
		                            "0110",
		                            "0111",
		                            "1000",
		                            "1001",
		                            "1010",
		                            "1011",
		                            "1100",
		                            "1101",
		                            "1110",
		                            "1111");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 27 :: 10 | 14 --
	end generate;
    gen_mcs_rom_27: if sel = 27 generate

		constant MEMORY : v_arr := ("0000",
		                            "1010",
		                            "0111",
		                            "1101",
		                            "1110",
		                            "0100",
		                            "1001",
		                            "0011",
		                            "1111",
		                            "0101",
		                            "1000",
		                            "0010",
		                            "0001",
		                            "1011",
		                            "0110",
		                            "1100",
		                            "0000",
		                            "1110",
		                            "1111",
		                            "0001",
		                            "1101",
		                            "0011",
		                            "0010",
		                            "1100",
		                            "1001",
		                            "0111",
		                            "0110",
		                            "1000",
		                            "0100",
		                            "1010",
		                            "1011",
		                            "0101");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 28 :: 15 | 5 --
	end generate;
    gen_mcs_rom_28: if sel = 28 generate

		constant MEMORY : v_arr := ("0000",
		                            "1111",
		                            "1101",
		                            "0010",
		                            "1001",
		                            "0110",
		                            "0100",
		                            "1011",
		                            "0001",
		                            "1110",
		                            "1100",
		                            "0011",
		                            "1000",
		                            "0111",
		                            "0101",
		                            "1010",
		                            "0000",
		                            "0101",
		                            "1010",
		                            "1111",
		                            "0111",
		                            "0010",
		                            "1101",
		                            "1000",
		                            "1110",
		                            "1011",
		                            "0100",
		                            "0001",
		                            "1001",
		                            "1100",
		                            "0011",
		                            "0110");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 29 :: 1 | 10 --
	end generate;
    gen_mcs_rom_29: if sel = 29 generate

		constant MEMORY : v_arr := ("0000",
		                            "0001",
		                            "0010",
		                            "0011",
		                            "0100",
		                            "0101",
		                            "0110",
		                            "0111",
		                            "1000",
		                            "1001",
		                            "1010",
		                            "1011",
		                            "1100",
		                            "1101",
		                            "1110",
		                            "1111",
		                            "0000",
		                            "1010",
		                            "0111",
		                            "1101",
		                            "1110",
		                            "0100",
		                            "1001",
		                            "0011",
		                            "1111",
		                            "0101",
		                            "1000",
		                            "0010",
		                            "0001",
		                            "1011",
		                            "0110",
		                            "1100");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 30 :: 13 | 2 --
	end generate;
    gen_mcs_rom_30: if sel = 30 generate

		constant MEMORY : v_arr := ("0000",
		                            "1101",
		                            "1001",
		                            "0100",
		                            "0001",
		                            "1100",
		                            "1000",
		                            "0101",
		                            "0010",
		                            "1111",
		                            "1011",
		                            "0110",
		                            "0011",
		                            "1110",
		                            "1010",
		                            "0111",
		                            "0000",
		                            "0010",
		                            "0100",
		                            "0110",
		                            "1000",
		                            "1010",
		                            "1100",
		                            "1110",
		                            "0011",
		                            "0001",
		                            "0111",
		                            "0101",
		                            "1011",
		                            "1001",
		                            "1111",
		                            "1101");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);

	-- Cell 31 :: 10 | 3 --
	end generate;
    gen_mcs_rom_31: if sel = 31 generate

		constant MEMORY : v_arr := ("0000",
		                            "1010",
		                            "0111",
		                            "1101",
		                            "1110",
		                            "0100",
		                            "1001",
		                            "0011",
		                            "1111",
		                            "0101",
		                            "1000",
		                            "0010",
		                            "0001",
		                            "1011",
		                            "0110",
		                            "1100",
		                            "0000",
		                            "0011",
		                            "0110",
		                            "0101",
		                            "1100",
		                            "1111",
		                            "1010",
		                            "1001",
		                            "1011",
		                            "1000",
		                            "1101",
		                            "1110",
		                            "0111",
		                            "0100",
		                            "0001",
		                            "0010");

	begin
		input1 <= to_integer(unsigned(ADDR));
		Dout   <= MEMORY(input1);
	end generate;
end mr0;
